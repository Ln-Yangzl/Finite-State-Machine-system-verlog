`ifndef __LAB6_SVH
`define __LAB6_SVH

typedef enum logic [1:0] {
     GREEN_RED, YELLOW_RED, RED_GREEN, RED_YELLOW 
} state_t;

`endif
